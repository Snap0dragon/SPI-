interface spi_if;
  logic mosi;  
  logic miso;  
  logic sclk; 
  logic cs;    
endinterface